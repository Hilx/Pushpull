LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

PACKAGE dsl_pack_func IS
  FUNCTION MAXIMUM(X, Y : INTEGER) RETURN INTEGER;
END PACKAGE;

PACKAGE BODY dsl_pack_func IS
  
  FUNCTION MAXIMUM(X, Y : INTEGER) RETURN INTEGER IS
    VARIABLE Z : INTEGER;
  BEGIN
    IF X > Y THEN
      Z := X;
    ELSE
      Z := Y;
    END IF;
    RETURN Z;
  END FUNCTION;
  
END PACKAGE BODY;
